<svg width="30" height="22" viewBox="0 0 30 22" fill="none" xmlns="http://www.w3.org/2000/svg">
<path d="M29.9294 16.7188C29.93 16.7129 29.93 16.7071 29.9294 16.7013L27.8806 6.18C27.8806 6.1725 27.8806 6.165 27.8806 6.1575C27.5644 4.43007 26.6527 2.86809 25.3042 1.74314C23.9556 0.618184 22.2555 0.00139391 20.4994 5.53315e-07H9.48562C7.72455 -0.000676284 6.01964 0.619617 4.67073 1.75179C3.32182 2.88395 2.41531 4.45549 2.11062 6.19L0.0718687 16.7013C0.0712666 16.7071 0.0712666 16.7129 0.0718687 16.7188C-0.0940781 17.661 0.0446289 18.6317 0.467851 19.4898C0.891073 20.3479 1.57678 21.0487 2.42541 21.4906C3.27405 21.9325 4.24143 22.0924 5.18711 21.947C6.1328 21.8017 7.00755 21.3588 7.68437 20.6825L7.72812 20.6362L12.6894 15H17.3144L22.2781 20.6362C22.2919 20.6525 22.3069 20.6675 22.3219 20.6825C23.1654 21.5242 24.3077 21.9979 25.4994 22C26.1562 21.9996 26.805 21.8554 27.4002 21.5775C27.9954 21.2996 28.5225 20.8948 28.9445 20.3915C29.3666 19.8882 29.6734 19.2986 29.8433 18.6641C30.0132 18.0296 30.0422 17.3656 29.9281 16.7188H29.9294ZM11.9994 9H10.9994V10C10.9994 10.2652 10.894 10.5196 10.7065 10.7071C10.5189 10.8946 10.2646 11 9.99937 11C9.73415 11 9.4798 10.8946 9.29226 10.7071C9.10473 10.5196 8.99937 10.2652 8.99937 10V9H7.99937C7.73415 9 7.4798 8.89464 7.29226 8.70711C7.10473 8.51957 6.99937 8.26522 6.99937 8C6.99937 7.73478 7.10473 7.48043 7.29226 7.29289C7.4798 7.10536 7.73415 7 7.99937 7H8.99937V6C8.99937 5.73478 9.10473 5.48043 9.29226 5.29289C9.4798 5.10536 9.73415 5 9.99937 5C10.2646 5 10.5189 5.10536 10.7065 5.29289C10.894 5.48043 10.9994 5.73478 10.9994 6V7H11.9994C12.2646 7 12.5189 7.10536 12.7065 7.29289C12.894 7.48043 12.9994 7.73478 12.9994 8C12.9994 8.26522 12.894 8.51957 12.7065 8.70711C12.5189 8.89464 12.2646 9 11.9994 9ZM16.9994 8C16.9994 7.73478 17.1047 7.48043 17.2923 7.29289C17.4798 7.10536 17.7342 7 17.9994 7H20.9994C21.2646 7 21.5189 7.10536 21.7065 7.29289C21.894 7.48043 21.9994 7.73478 21.9994 8C21.9994 8.26522 21.894 8.51957 21.7065 8.70711C21.5189 8.89464 21.2646 9 20.9994 9H17.9994C17.7342 9 17.4798 8.89464 17.2923 8.70711C17.1047 8.51957 16.9994 8.26522 16.9994 8ZM27.5456 18.9338C27.3583 19.2034 27.1193 19.4332 26.8425 19.6098C26.5657 19.7864 26.2566 19.9063 25.9331 19.9625C25.5418 20.0309 25.1398 20.0056 24.7602 19.8884C24.3805 19.7713 24.0341 19.5658 23.7494 19.2887L19.9744 15H20.4994C21.7761 15.0002 23.0317 14.6744 24.1473 14.0536C25.2629 13.4328 26.2015 12.5375 26.8744 11.4525L27.9669 17.0775C28.0225 17.3994 28.0139 17.7291 27.9416 18.0477C27.8693 18.3663 27.7347 18.6674 27.5456 18.9338Z" fill="url(#paint0_linear_2213_669)"/>



<defs>
<linearGradient id="paint0_linear_2213_669" x1="0.00366211" y1="11" x2="29.9965" y2="11" gradientUnits="userSpaceOnUse">
<stop stop-color="#FC4A1A"/>
<stop offset="1" stop-color="#F7B733"/>
</linearGradient>
</defs>
</svg>
